magic
tech scmos
timestamp 1612710923
<< nwell >>
rect -36 11 -15 15
rect -36 -6 17 11
rect -36 -9 -15 -6
<< ntransistor >>
rect -25 26 -22 28
rect -4 17 -2 20
rect 4 17 6 20
<< ptransistor >>
rect -24 2 -21 4
rect -4 2 -2 5
rect 4 2 6 5
<< ndiffusion >>
rect -25 28 -22 29
rect -25 25 -22 26
rect -5 17 -4 20
rect -2 17 -1 20
rect 3 17 4 20
rect 6 17 7 20
<< pdiffusion >>
rect -24 4 -21 5
rect -24 1 -21 2
rect -5 2 -4 5
rect -2 2 -1 5
rect 3 2 4 5
rect 6 2 7 5
<< ndcontact >>
rect -26 29 -22 33
rect -26 21 -22 25
rect -9 17 -5 21
rect -1 17 3 21
rect 7 17 11 21
<< pdcontact >>
rect -25 5 -21 9
rect -9 1 -5 5
rect -25 -3 -21 1
rect -1 1 3 5
rect 7 1 11 5
<< psubstratepcontact >>
rect -5 25 -1 29
<< nsubstratencontact >>
rect -33 4 -29 8
<< polysilicon >>
rect -30 26 -25 28
rect -22 26 -18 28
rect -20 4 -18 26
rect -4 20 -2 22
rect 4 20 6 22
rect -4 5 -2 17
rect 4 5 6 17
rect -26 2 -24 4
rect -21 2 -18 4
rect -4 -2 -2 2
rect 4 -2 6 2
<< polycontact >>
rect -18 1 -14 5
rect -5 -6 -1 -2
rect 3 -6 7 -2
<< metal1 >>
rect -1 29 3 33
rect -25 9 -22 17
rect -18 18 -9 21
rect -18 14 -15 18
rect -18 11 3 14
rect -18 5 -15 11
rect 0 5 3 11
rect -32 -2 -29 4
rect -10 4 -9 5
rect -11 1 -9 4
rect -11 -2 -8 1
<< m2contact >>
rect -22 29 -18 33
rect -1 25 3 29
rect 7 21 11 25
rect -26 17 -22 21
rect 7 5 11 9
rect -29 -3 -25 1
rect -12 -6 -8 -2
rect -5 -10 -1 -6
rect 3 -10 7 -6
<< metal2 >>
rect -18 28 -15 32
rect -18 25 -1 28
rect 3 25 10 28
rect -29 5 7 8
rect -29 1 -26 5
rect -12 -2 -9 5
<< m3contact >>
rect -30 17 -26 21
rect -5 -14 -1 -10
rect 4 -14 8 -10
<< metal3 >>
rect -31 21 -25 22
rect -31 17 -30 21
rect -26 17 -25 21
rect -31 16 -25 17
rect -6 -10 0 -9
rect -6 -14 -5 -10
rect -1 -14 0 -10
rect -6 -15 0 -14
rect 3 -10 9 -9
rect 3 -14 4 -10
rect 8 -14 9 -10
rect 3 -15 9 -14
<< labels >>
rlabel m3contact -28 19 -28 19 1 out
rlabel metal1 -31 1 -31 1 3 Vdd
rlabel metal1 1 31 1 31 5 Gnd
rlabel m3contact -3 -12 -3 -12 1 in1
rlabel m3contact 5 -12 5 -12 1 in2
<< end >>
