magic
tech scmos
timestamp 1605897077
<< nwell >>
rect -7 11 12 40
<< ntransistor >>
rect 0 -2 6 0
<< ptransistor >>
rect 0 22 6 24
<< ndiffusion >>
rect 0 1 1 4
rect 5 1 6 4
rect 0 0 6 1
rect 0 -3 6 -2
rect 0 -6 1 -3
rect 5 -6 6 -3
<< pdiffusion >>
rect 0 25 1 28
rect 5 25 6 28
rect 0 24 6 25
rect 0 21 6 22
rect 0 18 1 21
rect 5 18 6 21
<< ndcontact >>
rect 1 1 5 5
rect 1 -7 5 -3
<< pdcontact >>
rect 1 25 5 29
rect 1 17 5 21
<< psubstratepcontact >>
rect 1 -15 5 -11
<< nsubstratencontact >>
rect 1 33 5 37
<< polysilicon >>
rect -2 22 0 24
rect 6 22 8 24
rect -2 -2 0 0
rect 6 -2 8 0
<< polycontact >>
rect -6 21 -2 25
rect -6 -3 -2 1
<< metal1 >>
rect -7 33 1 37
rect 5 33 12 37
rect -7 32 12 33
rect 1 29 5 32
rect -6 1 -3 21
rect 2 12 5 17
rect 2 9 12 12
rect 2 5 5 9
rect 1 -10 5 -7
rect -7 -11 12 -10
rect -7 -15 1 -11
rect 5 -15 12 -11
<< labels >>
rlabel metal1 -5 10 -5 10 1 in
rlabel metal1 8 10 8 10 1 out
rlabel metal1 -5 -13 -5 -13 2 Gnd
rlabel metal1 -5 34 -5 34 3 Vdd
<< end >>
