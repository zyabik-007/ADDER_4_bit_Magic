* Podstawowy test sumatora 4-bitowego - test dodawania A+B=S przy 1 MHz.
* Test wykonuje dodawania 0000+0000 oraz 1111+1111 naprzemiennie co 0.5 us.

.lib .\scn05mos59_ltspice.lib

.include ADDER4bit.spice

Vdd vdd 0 dc 3
Vshort gnd 0 dc 0

** dodatkowe obciazenie wyjsc
.subckt INV in out vdd
  M1 out in 0 0 nfet w=1.8u l=0.6u
  M2 out in vdd vdd pfet w=1.8u l=0.6u
.ends

x10 S0 S0_ vdd INV
x20 S1 S1_ vdd INV
x30 S2 S2_ vdd INV
x40 S3 S3_ vdd INV
x50 S4 S4_ vdd INV

************************

VA0 A0 0 dc 0 pulse(0 3 0.5u 1n 1n 0.5u 1u)
VA1 A1 0 dc 0 pulse(0 3 0.5u 1n 1n 0.5u 1u)
VA2 A2 0 dc 0 pulse(0 3 0.5u 1n 1n 0.5u 1u)
VA3 A3 0 dc 0 pulse(0 3 0.5u 1n 1n 0.5u 1u)

VB0 B0 0 dc 0 pulse(0 3 0.5u 1n 1n 0.5u 1u)
VB1 B1 0 dc 0 pulse(0 3 0.5u 1n 1n 0.5u 1u)
VB2 B2 0 dc 0 pulse(0 3 0.5u 1n 1n 0.5u 1u)
VB3 B3 0 dc 0 pulse(0 3 0.5u 1n 1n 0.5u 1u)

.op
.tran 1u 2u 0
.probe v([S0]) v([S1]) v([S2]) v([S3]) v([S4])
.end


