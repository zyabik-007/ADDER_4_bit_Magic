* Test szybkosci sumatora 4-bitowego - test dodawania A+B=S przy 1000 MHz
* Test wykonuje dodawania 0000+0000 oraz 1111+1111 naprzemiennie co 1/2 ns

.lib .\scn05mos59_ltspice.lib

.include ADDER4bit.spice

Vdd vdd 0 dc 3
Vshort gnd 0 dc 0

** Dodatkowe obciazenie wyjsc *************

.subckt INV in out vdd
  M1 out in 0 0 nfet w=1.8u l=0.6u
  M2 out in vdd vdd pfet w=1.8u l=0.6u
.ends

.subckt XOR2 in1 in2 out vdd
M1 out in2 1   0     NFET W=1.8u L=0.6u
M2 out in2 in1 vdd   PFET W=1.8u L=0.6u
M3 out 1   in2 0     NFET W=1.8u L=0.6u
M4 out in1 in2 vdd   PFET W=1.8u L=0.6u
M5 1   in1 0   0     NFET W=1.8u L=0.6u
M6 1   in1 vdd vdd   PFET W=1.8u L=0.6u
.ends

.subckt OR2 in1 in2 out vdd
M1 1   in1 vdd vdd   PFET W=1.8u L=0.6u
M2 2   in2 1   vdd   PFET W=1.8u L=0.6u
M3 2   in1 0   0     NFET W=1.8u L=0.6u
M4 2   in2 0   0     NFET W=1.8u L=0.6u
M5 out 2   vdd vdd   PFET W=1.8u L=0.6u
M6 out 2   0   0     NFET W=1.8u L=0.6u
.ends

.subckt AND2 in1 in2 out vdd
M1 1   in1 vdd vdd   PFET W=1.8u L=0.6u
M2 1   in2 vdd vdd   PFET W=1.8u L=0.6u
M3 1   in1 2   0     NFET W=1.8u L=0.6u
M4 2   in2 0   0     NFET W=1.8u L=0.6u
M5 out 1   vdd vdd   PFET W=1.8u L=0.6u
M6 out 1   0   0     NFET W=1.8u L=0.6u
.ends


.subckt ADDER1bit in1 in2 Cin out Cout vdd
x1 in1 in2  1    vdd   xor2
x2 1   Cin  out  vdd   xor2
x3 1   Cin  2    vdd   and2
x4 in1 in2  3    vdd   and2
x5 2   3    Cout vdd   or2
.ends


x10 S0 S0_ vdd INV
x20 S1 S1_ vdd INV
x30 S2 S2_ vdd INV
x40 S3 S3_ vdd INV
x50 S4 S4_ vdd INV
x55 0 0 S4 out_ Cout_ vdd ADDER1bit
***Koniec: dodatkowe obciazenie wyjsc*********************

.param period=1ns

VA A 0 dc 0 pulse(0 3 {period/2} {period/50} {period/50} {period/2} {period})
RA0 A0 A 1
RA1 A1 A 1
RA2 A2 A 1
RA3 A3 A 1

VB B 0 dc 0 pulse(0 3 {period/2} {period/50} {period/50} {period/2} {period})
RB0 B0 B 1
RB1 B1 B 1
RB2 B2 B 1
RB3 B3 B 1


.op
.tran 1n 4n 0
.probe v([S4]) v([A]) v([B])
.end


